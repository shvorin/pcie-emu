// pcie_de_gen1_x8_ast128.v

// Generated using ACDS version 12.1 177 at 2013.02.08.15:37:13

`timescale 1 ps / 1 ps
module pcie_de_gen1_x8_ast128 (
		input  wire        refclk_clk,                //     refclk.clk
		input  wire [31:0] hip_ctrl_test_in,          //   hip_ctrl.test_in
		input  wire        hip_ctrl_simu_mode_pipe,   //           .simu_mode_pipe
		input  wire        hip_serial_rx_in0,         // hip_serial.rx_in0
		input  wire        hip_serial_rx_in1,         //           .rx_in1
		input  wire        hip_serial_rx_in2,         //           .rx_in2
		input  wire        hip_serial_rx_in3,         //           .rx_in3
		input  wire        hip_serial_rx_in4,         //           .rx_in4
		input  wire        hip_serial_rx_in5,         //           .rx_in5
		input  wire        hip_serial_rx_in6,         //           .rx_in6
		input  wire        hip_serial_rx_in7,         //           .rx_in7
		output wire        hip_serial_tx_out0,        //           .tx_out0
		output wire        hip_serial_tx_out1,        //           .tx_out1
		output wire        hip_serial_tx_out2,        //           .tx_out2
		output wire        hip_serial_tx_out3,        //           .tx_out3
		output wire        hip_serial_tx_out4,        //           .tx_out4
		output wire        hip_serial_tx_out5,        //           .tx_out5
		output wire        hip_serial_tx_out6,        //           .tx_out6
		output wire        hip_serial_tx_out7,        //           .tx_out7
		input  wire        hip_pipe_sim_pipe_pclk_in, //   hip_pipe.sim_pipe_pclk_in
		output wire [1:0]  hip_pipe_sim_pipe_rate,    //           .sim_pipe_rate
		output wire [4:0]  hip_pipe_sim_ltssmstate,   //           .sim_ltssmstate
		output wire [2:0]  hip_pipe_eidleinfersel0,   //           .eidleinfersel0
		output wire [2:0]  hip_pipe_eidleinfersel1,   //           .eidleinfersel1
		output wire [2:0]  hip_pipe_eidleinfersel2,   //           .eidleinfersel2
		output wire [2:0]  hip_pipe_eidleinfersel3,   //           .eidleinfersel3
		output wire [2:0]  hip_pipe_eidleinfersel4,   //           .eidleinfersel4
		output wire [2:0]  hip_pipe_eidleinfersel5,   //           .eidleinfersel5
		output wire [2:0]  hip_pipe_eidleinfersel6,   //           .eidleinfersel6
		output wire [2:0]  hip_pipe_eidleinfersel7,   //           .eidleinfersel7
		output wire [1:0]  hip_pipe_powerdown0,       //           .powerdown0
		output wire [1:0]  hip_pipe_powerdown1,       //           .powerdown1
		output wire [1:0]  hip_pipe_powerdown2,       //           .powerdown2
		output wire [1:0]  hip_pipe_powerdown3,       //           .powerdown3
		output wire [1:0]  hip_pipe_powerdown4,       //           .powerdown4
		output wire [1:0]  hip_pipe_powerdown5,       //           .powerdown5
		output wire [1:0]  hip_pipe_powerdown6,       //           .powerdown6
		output wire [1:0]  hip_pipe_powerdown7,       //           .powerdown7
		output wire        hip_pipe_rxpolarity0,      //           .rxpolarity0
		output wire        hip_pipe_rxpolarity1,      //           .rxpolarity1
		output wire        hip_pipe_rxpolarity2,      //           .rxpolarity2
		output wire        hip_pipe_rxpolarity3,      //           .rxpolarity3
		output wire        hip_pipe_rxpolarity4,      //           .rxpolarity4
		output wire        hip_pipe_rxpolarity5,      //           .rxpolarity5
		output wire        hip_pipe_rxpolarity6,      //           .rxpolarity6
		output wire        hip_pipe_rxpolarity7,      //           .rxpolarity7
		output wire        hip_pipe_txcompl0,         //           .txcompl0
		output wire        hip_pipe_txcompl1,         //           .txcompl1
		output wire        hip_pipe_txcompl2,         //           .txcompl2
		output wire        hip_pipe_txcompl3,         //           .txcompl3
		output wire        hip_pipe_txcompl4,         //           .txcompl4
		output wire        hip_pipe_txcompl5,         //           .txcompl5
		output wire        hip_pipe_txcompl6,         //           .txcompl6
		output wire        hip_pipe_txcompl7,         //           .txcompl7
		output wire [7:0]  hip_pipe_txdata0,          //           .txdata0
		output wire [7:0]  hip_pipe_txdata1,          //           .txdata1
		output wire [7:0]  hip_pipe_txdata2,          //           .txdata2
		output wire [7:0]  hip_pipe_txdata3,          //           .txdata3
		output wire [7:0]  hip_pipe_txdata4,          //           .txdata4
		output wire [7:0]  hip_pipe_txdata5,          //           .txdata5
		output wire [7:0]  hip_pipe_txdata6,          //           .txdata6
		output wire [7:0]  hip_pipe_txdata7,          //           .txdata7
		output wire        hip_pipe_txdatak0,         //           .txdatak0
		output wire        hip_pipe_txdatak1,         //           .txdatak1
		output wire        hip_pipe_txdatak2,         //           .txdatak2
		output wire        hip_pipe_txdatak3,         //           .txdatak3
		output wire        hip_pipe_txdatak4,         //           .txdatak4
		output wire        hip_pipe_txdatak5,         //           .txdatak5
		output wire        hip_pipe_txdatak6,         //           .txdatak6
		output wire        hip_pipe_txdatak7,         //           .txdatak7
		output wire        hip_pipe_txdetectrx0,      //           .txdetectrx0
		output wire        hip_pipe_txdetectrx1,      //           .txdetectrx1
		output wire        hip_pipe_txdetectrx2,      //           .txdetectrx2
		output wire        hip_pipe_txdetectrx3,      //           .txdetectrx3
		output wire        hip_pipe_txdetectrx4,      //           .txdetectrx4
		output wire        hip_pipe_txdetectrx5,      //           .txdetectrx5
		output wire        hip_pipe_txdetectrx6,      //           .txdetectrx6
		output wire        hip_pipe_txdetectrx7,      //           .txdetectrx7
		output wire        hip_pipe_txelecidle0,      //           .txelecidle0
		output wire        hip_pipe_txelecidle1,      //           .txelecidle1
		output wire        hip_pipe_txelecidle2,      //           .txelecidle2
		output wire        hip_pipe_txelecidle3,      //           .txelecidle3
		output wire        hip_pipe_txelecidle4,      //           .txelecidle4
		output wire        hip_pipe_txelecidle5,      //           .txelecidle5
		output wire        hip_pipe_txelecidle6,      //           .txelecidle6
		output wire        hip_pipe_txelecidle7,      //           .txelecidle7
		output wire        hip_pipe_txdeemph0,        //           .txdeemph0
		output wire        hip_pipe_txdeemph1,        //           .txdeemph1
		output wire        hip_pipe_txdeemph2,        //           .txdeemph2
		output wire        hip_pipe_txdeemph3,        //           .txdeemph3
		output wire        hip_pipe_txdeemph4,        //           .txdeemph4
		output wire        hip_pipe_txdeemph5,        //           .txdeemph5
		output wire        hip_pipe_txdeemph6,        //           .txdeemph6
		output wire        hip_pipe_txdeemph7,        //           .txdeemph7
		output wire [2:0]  hip_pipe_txmargin0,        //           .txmargin0
		output wire [2:0]  hip_pipe_txmargin1,        //           .txmargin1
		output wire [2:0]  hip_pipe_txmargin2,        //           .txmargin2
		output wire [2:0]  hip_pipe_txmargin3,        //           .txmargin3
		output wire [2:0]  hip_pipe_txmargin4,        //           .txmargin4
		output wire [2:0]  hip_pipe_txmargin5,        //           .txmargin5
		output wire [2:0]  hip_pipe_txmargin6,        //           .txmargin6
		output wire [2:0]  hip_pipe_txmargin7,        //           .txmargin7
		output wire        hip_pipe_txswing0,         //           .txswing0
		output wire        hip_pipe_txswing1,         //           .txswing1
		output wire        hip_pipe_txswing2,         //           .txswing2
		output wire        hip_pipe_txswing3,         //           .txswing3
		output wire        hip_pipe_txswing4,         //           .txswing4
		output wire        hip_pipe_txswing5,         //           .txswing5
		output wire        hip_pipe_txswing6,         //           .txswing6
		output wire        hip_pipe_txswing7,         //           .txswing7
		input  wire        hip_pipe_phystatus0,       //           .phystatus0
		input  wire        hip_pipe_phystatus1,       //           .phystatus1
		input  wire        hip_pipe_phystatus2,       //           .phystatus2
		input  wire        hip_pipe_phystatus3,       //           .phystatus3
		input  wire        hip_pipe_phystatus4,       //           .phystatus4
		input  wire        hip_pipe_phystatus5,       //           .phystatus5
		input  wire        hip_pipe_phystatus6,       //           .phystatus6
		input  wire        hip_pipe_phystatus7,       //           .phystatus7
		input  wire [7:0]  hip_pipe_rxdata0,          //           .rxdata0
		input  wire [7:0]  hip_pipe_rxdata1,          //           .rxdata1
		input  wire [7:0]  hip_pipe_rxdata2,          //           .rxdata2
		input  wire [7:0]  hip_pipe_rxdata3,          //           .rxdata3
		input  wire [7:0]  hip_pipe_rxdata4,          //           .rxdata4
		input  wire [7:0]  hip_pipe_rxdata5,          //           .rxdata5
		input  wire [7:0]  hip_pipe_rxdata6,          //           .rxdata6
		input  wire [7:0]  hip_pipe_rxdata7,          //           .rxdata7
		input  wire        hip_pipe_rxdatak0,         //           .rxdatak0
		input  wire        hip_pipe_rxdatak1,         //           .rxdatak1
		input  wire        hip_pipe_rxdatak2,         //           .rxdatak2
		input  wire        hip_pipe_rxdatak3,         //           .rxdatak3
		input  wire        hip_pipe_rxdatak4,         //           .rxdatak4
		input  wire        hip_pipe_rxdatak5,         //           .rxdatak5
		input  wire        hip_pipe_rxdatak6,         //           .rxdatak6
		input  wire        hip_pipe_rxdatak7,         //           .rxdatak7
		input  wire        hip_pipe_rxelecidle0,      //           .rxelecidle0
		input  wire        hip_pipe_rxelecidle1,      //           .rxelecidle1
		input  wire        hip_pipe_rxelecidle2,      //           .rxelecidle2
		input  wire        hip_pipe_rxelecidle3,      //           .rxelecidle3
		input  wire        hip_pipe_rxelecidle4,      //           .rxelecidle4
		input  wire        hip_pipe_rxelecidle5,      //           .rxelecidle5
		input  wire        hip_pipe_rxelecidle6,      //           .rxelecidle6
		input  wire        hip_pipe_rxelecidle7,      //           .rxelecidle7
		input  wire [2:0]  hip_pipe_rxstatus0,        //           .rxstatus0
		input  wire [2:0]  hip_pipe_rxstatus1,        //           .rxstatus1
		input  wire [2:0]  hip_pipe_rxstatus2,        //           .rxstatus2
		input  wire [2:0]  hip_pipe_rxstatus3,        //           .rxstatus3
		input  wire [2:0]  hip_pipe_rxstatus4,        //           .rxstatus4
		input  wire [2:0]  hip_pipe_rxstatus5,        //           .rxstatus5
		input  wire [2:0]  hip_pipe_rxstatus6,        //           .rxstatus6
		input  wire [2:0]  hip_pipe_rxstatus7,        //           .rxstatus7
		input  wire        hip_pipe_rxvalid0,         //           .rxvalid0
		input  wire        hip_pipe_rxvalid1,         //           .rxvalid1
		input  wire        hip_pipe_rxvalid2,         //           .rxvalid2
		input  wire        hip_pipe_rxvalid3,         //           .rxvalid3
		input  wire        hip_pipe_rxvalid4,         //           .rxvalid4
		input  wire        hip_pipe_rxvalid5,         //           .rxvalid5
		input  wire        hip_pipe_rxvalid6,         //           .rxvalid6
		input  wire        hip_pipe_rxvalid7,         //           .rxvalid7
		input  wire        pcie_rstn_npor,            //  pcie_rstn.npor
		input  wire        pcie_rstn_pin_perst,       //           .pin_perst
		input  wire        reset_reset_n,             //      reset.reset_n
		input  wire        clk_clk                    //        clk.clk
	);

	wire          apps_int_msi_app_msi_req;                              // APPS:app_msi_req -> DUT:app_msi_req
	wire          dut_int_msi_app_msi_ack;                               // DUT:app_msi_ack -> APPS:app_msi_ack
	wire    [0:0] apps_int_msi_app_int_sts;                              // APPS:app_int_sts -> DUT:app_int_sts
	wire          dut_int_msi_app_int_ack;                               // DUT:app_int_ack -> APPS:app_int_ack
	wire    [2:0] apps_int_msi_app_msi_tc;                               // APPS:app_msi_tc -> DUT:app_msi_tc
	wire    [4:0] apps_int_msi_app_msi_num;                              // APPS:app_msi_num -> DUT:app_msi_num
	wire          dut_hip_rst_serdes_pll_locked;                         // DUT:serdes_pll_locked -> APPS:serdes_pll_locked
	wire          apps_hip_rst_pld_core_ready;                           // APPS:pld_core_ready -> DUT:pld_core_ready
	wire          dut_hip_rst_pld_clk_inuse;                             // DUT:pld_clk_inuse -> APPS:pld_clk_inuse
	wire          dut_hip_rst_reset_status;                              // DUT:reset_status -> APPS:reset_status
	wire          dut_hip_rst_testin_zero;                               // DUT:testin_zero -> APPS:testin_zero
	wire          apps_config_tl_cpl_pending;                            // APPS:cpl_pending -> DUT:cpl_pending
	wire   [52:0] dut_config_tl_tl_cfg_sts;                              // DUT:tl_cfg_sts -> APPS:tl_cfg_sts
	wire   [31:0] dut_config_tl_tl_cfg_ctl;                              // DUT:tl_cfg_ctl -> APPS:tl_cfg_ctl
	wire    [3:0] dut_config_tl_tl_cfg_add;                              // DUT:tl_cfg_add -> APPS:tl_cfg_add
	wire    [4:0] apps_config_tl_hpg_ctrler;                             // APPS:hpg_ctrler -> DUT:hpg_ctrler
	wire    [6:0] apps_config_tl_cpl_err;                                // APPS:cpl_err -> DUT:cpl_err
	wire          dut_power_mngt_pme_to_sr;                              // DUT:pme_to_sr -> APPS:pme_to_sr
	wire          apps_power_mngt_pm_auxpwr;                             // APPS:pm_auxpwr -> DUT:pm_auxpwr
	wire    [9:0] apps_power_mngt_pm_data;                               // APPS:pm_data -> DUT:pm_data
	wire          apps_power_mngt_pme_to_cr;                             // APPS:pme_to_cr -> DUT:pme_to_cr
	wire          apps_power_mngt_pm_event;                              // APPS:pm_event -> DUT:pm_event
	wire          dut_hip_status_ev128ns;                                // DUT:ev128ns -> APPS:ev128ns
	wire    [3:0] dut_hip_status_int_status;                             // DUT:int_status -> APPS:int_status
	wire          dut_hip_status_ev1us;                                  // DUT:ev1us -> APPS:ev1us
	wire          dut_hip_status_derr_cor_ext_rcv;                       // DUT:derr_cor_ext_rcv -> APPS:derr_cor_ext_rcv
	wire    [4:0] dut_hip_status_ltssmstate;                             // DUT:ltssmstate -> APPS:ltssmstate
	wire          dut_hip_status_rx_par_err;                             // DUT:rx_par_err -> APPS:rx_par_err
	wire          dut_hip_status_derr_rpl;                               // DUT:derr_rpl -> APPS:derr_rpl
	wire          dut_hip_status_l2_exit;                                // DUT:l2_exit -> APPS:l2_exit
	wire          dut_hip_status_cfg_par_err;                            // DUT:cfg_par_err -> APPS:cfg_par_err
	wire    [3:0] dut_hip_status_lane_act;                               // DUT:lane_act -> APPS:lane_act
	wire          dut_hip_status_dlup_exit;                              // DUT:dlup_exit -> APPS:dlup_exit
	wire    [7:0] dut_hip_status_ko_cpl_spc_header;                      // DUT:ko_cpl_spc_header -> APPS:ko_cpl_spc_header
	wire          dut_hip_status_hotrst_exit;                            // DUT:hotrst_exit -> APPS:hotrst_exit
	wire   [11:0] dut_hip_status_ko_cpl_spc_data;                        // DUT:ko_cpl_spc_data -> APPS:ko_cpl_spc_data
	wire    [1:0] dut_hip_status_tx_par_err;                             // DUT:tx_par_err -> APPS:tx_par_err
	wire          dut_hip_status_dlup;                                   // DUT:dlup -> APPS:dlup
	wire          dut_hip_status_derr_cor_ext_rpl;                       // DUT:derr_cor_ext_rpl -> APPS:derr_cor_ext_rpl
	wire   [11:0] dut_tx_cred_tx_cred_datafccp;                          // DUT:tx_cred_datafccp -> APPS:tx_cred_datafccp
	wire    [7:0] dut_tx_cred_tx_cred_hdrfcnp;                           // DUT:tx_cred_hdrfcnp -> APPS:tx_cred_hdrfcnp
	wire    [7:0] dut_tx_cred_tx_cred_hdrfccp;                           // DUT:tx_cred_hdrfccp -> APPS:tx_cred_hdrfccp
	wire    [5:0] dut_tx_cred_tx_cred_fchipcons;                         // DUT:tx_cred_fchipcons -> APPS:tx_cred_fchipcons
	wire    [7:0] dut_tx_cred_tx_cred_hdrfcp;                            // DUT:tx_cred_hdrfcp -> APPS:tx_cred_hdrfcp
	wire   [11:0] dut_tx_cred_tx_cred_datafcp;                           // DUT:tx_cred_datafcp -> APPS:tx_cred_datafcp
	wire    [5:0] dut_tx_cred_tx_cred_fcinfinite;                        // DUT:tx_cred_fcinfinite -> APPS:tx_cred_fcinfinite
	wire   [11:0] dut_tx_cred_tx_cred_datafcnp;                          // DUT:tx_cred_datafcnp -> APPS:tx_cred_datafcnp
	wire          apps_rx_bar_be_rx_st_mask;                             // APPS:rx_st_mask -> DUT:rx_st_mask
	wire   [15:0] dut_rx_bar_be_rx_st_be;                                // DUT:rx_st_be -> APPS:rx_st_be
	wire    [7:0] dut_rx_bar_be_rx_st_bar;                               // DUT:rx_st_bar -> APPS:rx_st_bar
	wire    [0:0] apps_tx_st_endofpacket;                                // APPS:tx_st_eop -> DUT:tx_st_eop
	wire    [0:0] apps_tx_st_valid;                                      // APPS:tx_st_valid -> DUT:tx_st_valid
	wire    [0:0] apps_tx_st_startofpacket;                              // APPS:tx_st_sop -> DUT:tx_st_sop
	wire    [0:0] apps_tx_st_error;                                      // APPS:tx_st_err -> DUT:tx_st_err
	wire  [127:0] apps_tx_st_data;                                       // APPS:tx_st_data -> DUT:tx_st_data
	wire    [1:0] apps_tx_st_empty;                                      // APPS:tx_st_empty -> DUT:tx_st_empty
	wire          apps_tx_st_ready;                                      // DUT:tx_st_ready -> APPS:tx_st_ready
	wire   [31:0] dut_lmi_lmi_dout;                                      // DUT:lmi_dout -> APPS:lmi_dout
	wire          apps_lmi_lmi_wren;                                     // APPS:lmi_wren -> DUT:lmi_wren
	wire   [31:0] apps_lmi_lmi_din;                                      // APPS:lmi_din -> DUT:lmi_din
	wire          apps_lmi_lmi_rden;                                     // APPS:lmi_rden -> DUT:lmi_rden
	wire   [11:0] apps_lmi_lmi_addr;                                     // APPS:lmi_addr -> DUT:lmi_addr
	wire          dut_lmi_lmi_ack;                                       // DUT:lmi_ack -> APPS:lmi_ack
	wire    [0:0] dut_rx_st_endofpacket;                                 // DUT:rx_st_eop -> APPS:rx_st_eop
	wire    [0:0] dut_rx_st_valid;                                       // DUT:rx_st_valid -> APPS:rx_st_valid
	wire    [0:0] dut_rx_st_startofpacket;                               // DUT:rx_st_sop -> APPS:rx_st_sop
	wire    [0:0] dut_rx_st_error;                                       // DUT:rx_st_err -> APPS:rx_st_err
	wire  [127:0] dut_rx_st_data;                                        // DUT:rx_st_data -> APPS:rx_st_data
	wire    [1:0] dut_rx_st_empty;                                       // DUT:rx_st_empty -> APPS:rx_st_empty
	wire          dut_rx_st_ready;                                       // APPS:rx_st_ready -> DUT:rx_st_ready
	wire          apps_pld_clk_hip_clk;                                  // APPS:pld_clk_hip -> [DUT:pld_clk, pcie_reconfig_driver_0:pld_clk]
	wire          dut_coreclkout_hip_clk;                                // DUT:coreclkout_hip -> APPS:coreclkout_hip
	wire  [459:0] dut_reconfig_from_xcvr_reconfig_from_xcvr;             // DUT:reconfig_from_xcvr -> alt_xcvr_reconfig_0:reconfig_from_xcvr
	wire  [699:0] alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr; // alt_xcvr_reconfig_0:reconfig_to_xcvr -> DUT:reconfig_to_xcvr
	wire          pcie_reconfig_driver_0_reconfig_mgmt_waitrequest;      // alt_xcvr_reconfig_0:reconfig_mgmt_waitrequest -> pcie_reconfig_driver_0:reconfig_mgmt_waitrequest
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_writedata;        // pcie_reconfig_driver_0:reconfig_mgmt_writedata -> alt_xcvr_reconfig_0:reconfig_mgmt_writedata
	wire    [6:0] pcie_reconfig_driver_0_reconfig_mgmt_address;          // pcie_reconfig_driver_0:reconfig_mgmt_address -> alt_xcvr_reconfig_0:reconfig_mgmt_address
	wire          pcie_reconfig_driver_0_reconfig_mgmt_write;            // pcie_reconfig_driver_0:reconfig_mgmt_write -> alt_xcvr_reconfig_0:reconfig_mgmt_write
	wire          pcie_reconfig_driver_0_reconfig_mgmt_read;             // pcie_reconfig_driver_0:reconfig_mgmt_read -> alt_xcvr_reconfig_0:reconfig_mgmt_read
	wire   [31:0] pcie_reconfig_driver_0_reconfig_mgmt_readdata;         // alt_xcvr_reconfig_0:reconfig_mgmt_readdata -> pcie_reconfig_driver_0:reconfig_mgmt_readdata
	wire    [1:0] dut_hip_currentspeed_currentspeed;                     // DUT:currentspeed -> pcie_reconfig_driver_0:currentspeed
	wire          alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy;       // alt_xcvr_reconfig_0:reconfig_busy -> pcie_reconfig_driver_0:reconfig_busy
	wire          apps_hip_status_drv_derr_rpl_drv;                      // APPS:derr_rpl_drv -> pcie_reconfig_driver_0:derr_rpl_drv
	wire    [4:0] apps_hip_status_drv_ltssmstate_drv;                    // APPS:ltssmstate_drv -> pcie_reconfig_driver_0:ltssmstate_drv
	wire          apps_hip_status_drv_dlup_exit_drv;                     // APPS:dlup_exit_drv -> pcie_reconfig_driver_0:dlup_exit_drv
	wire          apps_hip_status_drv_derr_cor_ext_rpl_drv;              // APPS:derr_cor_ext_rpl_drv -> pcie_reconfig_driver_0:derr_cor_ext_rpl_drv
	wire          apps_hip_status_drv_derr_cor_ext_rcv_drv;              // APPS:derr_cor_ext_rcv_drv -> pcie_reconfig_driver_0:derr_cor_ext_rcv_drv
	wire          apps_hip_status_drv_ev1us_drv;                         // APPS:ev1us_drv -> pcie_reconfig_driver_0:ev1us_drv
	wire    [3:0] apps_hip_status_drv_lane_act_drv;                      // APPS:lane_act_drv -> pcie_reconfig_driver_0:lane_act_drv
	wire          apps_hip_status_drv_l2_exit_drv;                       // APPS:l2_exit_drv -> pcie_reconfig_driver_0:l2_exit_drv
	wire    [3:0] apps_hip_status_drv_int_status_drv;                    // APPS:int_status_drv -> pcie_reconfig_driver_0:int_status_drv
	wire          apps_hip_status_drv_hotrst_exit_drv;                   // APPS:hotrst_exit_drv -> pcie_reconfig_driver_0:hotrst_exit_drv
	wire          apps_hip_status_drv_ev128ns_drv;                       // APPS:ev128ns_drv -> pcie_reconfig_driver_0:ev128ns_drv
	wire          rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [alt_xcvr_reconfig_0:mgmt_rst_reset, pcie_reconfig_driver_0:reconfig_xcvr_rst]

	altpcie_sv_hip_ast_hwtcl #(
		.lane_mask_hwtcl                          ("x8"),
		.gen123_lane_rate_mode_hwtcl              ("Gen1 (2.5 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.ast_width_hwtcl                          ("Avalon-ST 128-bit"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.use_ast_parity                           (0),
		.multiple_packets_per_cycle_hwtcl         (0),
		.in_cvp_mode_hwtcl                        (0),
		.use_pci_ext_hwtcl                        (0),
		.use_pcie_ext_hwtcl                       (0),
		.use_config_bypass_hwtcl                  (0),
		.hip_reconfig_hwtcl                       (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.bar0_size_mask_hwtcl                     (28),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Enabled"),
		.bar0_prefetchable_hwtcl                  ("Enabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (10),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.expansion_base_address_register_hwtcl    (0),
		.io_window_addr_width_hwtcl               (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.vendor_id_hwtcl                          (19283),
		.device_id_hwtcl                          (57345),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (3997696),
		.subsystem_vendor_id_hwtcl                (19283),
		.subsystem_device_id_hwtcl                (57345),
		.max_payload_size_hwtcl                   (256),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.rx_ei_l0s_hwtcl                          (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (40960),
		.vsec_rev_hwtcl                           (0),
		.reconfig_to_xcvr_width                   (700),
		.hip_hard_reset_hwtcl                     (1),
		.reconfig_from_xcvr_width                 (460),
		.single_rx_detect_hwtcl                   (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.sameclock_nfts_count_hwtcl               (128),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("true"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.aspm_config_management_hwtcl             ("true"),
		.millisecond_cycle_count_hwtcl            (124250),
		.deemphasis_enable_hwtcl                  ("false"),
		.port_width_be_hwtcl                      (16),
		.port_width_data_hwtcl                    (128),
		.gen3_dcbal_en_hwtcl                      (1),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.enable_pipe32_sim_hwtcl                  (0),
		.fixed_preset_on                          (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.bypass_clk_switch_hwtcl                  ("TRUE"),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.indicator_hwtcl                          (0),
		.enable_l1_aspm_hwtcl                     ("false"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.diffclock_nfts_count_hwtcl               (128),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.l2_async_logic_hwtcl                     ("disable"),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("true"),
		.atomic_malformed_hwtcl                   ("false"),
		.flr_capability_hwtcl                     ("true"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (195),
		.cpl_spc_data_hwtcl                       (781),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.hwtcl_override_g2_txvod                  (0),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15),
		.hwtcl_override_g3rxcoef                  (0),
		.gen3_coeff_1_hwtcl                       (7),
		.gen3_coeff_1_sel_hwtcl                   ("preset_1"),
		.gen3_coeff_1_preset_hint_hwtcl           (0),
		.gen3_coeff_1_nxtber_more_ptr_hwtcl       (1),
		.gen3_coeff_1_nxtber_more_hwtcl           ("g3_coeff_1_nxtber_more"),
		.gen3_coeff_1_nxtber_less_ptr_hwtcl       (1),
		.gen3_coeff_1_nxtber_less_hwtcl           ("g3_coeff_1_nxtber_less"),
		.gen3_coeff_1_reqber_hwtcl                (0),
		.gen3_coeff_1_ber_meas_hwtcl              (2),
		.gen3_coeff_2_hwtcl                       (0),
		.gen3_coeff_2_sel_hwtcl                   ("preset_2"),
		.gen3_coeff_2_preset_hint_hwtcl           (0),
		.gen3_coeff_2_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_2_nxtber_more_hwtcl           ("g3_coeff_2_nxtber_more"),
		.gen3_coeff_2_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_2_nxtber_less_hwtcl           ("g3_coeff_2_nxtber_less"),
		.gen3_coeff_2_reqber_hwtcl                (0),
		.gen3_coeff_2_ber_meas_hwtcl              (0),
		.gen3_coeff_3_hwtcl                       (0),
		.gen3_coeff_3_sel_hwtcl                   ("preset_3"),
		.gen3_coeff_3_preset_hint_hwtcl           (0),
		.gen3_coeff_3_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_3_nxtber_more_hwtcl           ("g3_coeff_3_nxtber_more"),
		.gen3_coeff_3_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_3_nxtber_less_hwtcl           ("g3_coeff_3_nxtber_less"),
		.gen3_coeff_3_reqber_hwtcl                (0),
		.gen3_coeff_3_ber_meas_hwtcl              (0),
		.gen3_coeff_4_hwtcl                       (0),
		.gen3_coeff_4_sel_hwtcl                   ("preset_4"),
		.gen3_coeff_4_preset_hint_hwtcl           (0),
		.gen3_coeff_4_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_4_nxtber_more_hwtcl           ("g3_coeff_4_nxtber_more"),
		.gen3_coeff_4_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_4_nxtber_less_hwtcl           ("g3_coeff_4_nxtber_less"),
		.gen3_coeff_4_reqber_hwtcl                (0),
		.gen3_coeff_4_ber_meas_hwtcl              (0),
		.gen3_coeff_5_hwtcl                       (0),
		.gen3_coeff_5_sel_hwtcl                   ("preset_5"),
		.gen3_coeff_5_preset_hint_hwtcl           (0),
		.gen3_coeff_5_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_5_nxtber_more_hwtcl           ("g3_coeff_5_nxtber_more"),
		.gen3_coeff_5_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_5_nxtber_less_hwtcl           ("g3_coeff_5_nxtber_less"),
		.gen3_coeff_5_reqber_hwtcl                (0),
		.gen3_coeff_5_ber_meas_hwtcl              (0),
		.gen3_coeff_6_hwtcl                       (0),
		.gen3_coeff_6_sel_hwtcl                   ("preset_6"),
		.gen3_coeff_6_preset_hint_hwtcl           (0),
		.gen3_coeff_6_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_6_nxtber_more_hwtcl           ("g3_coeff_6_nxtber_more"),
		.gen3_coeff_6_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_6_nxtber_less_hwtcl           ("g3_coeff_6_nxtber_less"),
		.gen3_coeff_6_reqber_hwtcl                (0),
		.gen3_coeff_6_ber_meas_hwtcl              (0),
		.gen3_coeff_7_hwtcl                       (0),
		.gen3_coeff_7_sel_hwtcl                   ("preset_7"),
		.gen3_coeff_7_preset_hint_hwtcl           (0),
		.gen3_coeff_7_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_7_nxtber_more_hwtcl           ("g3_coeff_7_nxtber_more"),
		.gen3_coeff_7_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_7_nxtber_less_hwtcl           ("g3_coeff_7_nxtber_less"),
		.gen3_coeff_7_reqber_hwtcl                (0),
		.gen3_coeff_7_ber_meas_hwtcl              (0),
		.gen3_coeff_8_hwtcl                       (0),
		.gen3_coeff_8_sel_hwtcl                   ("preset_8"),
		.gen3_coeff_8_preset_hint_hwtcl           (0),
		.gen3_coeff_8_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_8_nxtber_more_hwtcl           ("g3_coeff_8_nxtber_more"),
		.gen3_coeff_8_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_8_nxtber_less_hwtcl           ("g3_coeff_8_nxtber_less"),
		.gen3_coeff_8_reqber_hwtcl                (0),
		.gen3_coeff_8_ber_meas_hwtcl              (0),
		.gen3_coeff_9_hwtcl                       (0),
		.gen3_coeff_9_sel_hwtcl                   ("preset_9"),
		.gen3_coeff_9_preset_hint_hwtcl           (0),
		.gen3_coeff_9_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_9_nxtber_more_hwtcl           ("g3_coeff_9_nxtber_more"),
		.gen3_coeff_9_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_9_nxtber_less_hwtcl           ("g3_coeff_9_nxtber_less"),
		.gen3_coeff_9_reqber_hwtcl                (0),
		.gen3_coeff_9_ber_meas_hwtcl              (0),
		.gen3_coeff_10_hwtcl                      (0),
		.gen3_coeff_10_sel_hwtcl                  ("preset_10"),
		.gen3_coeff_10_preset_hint_hwtcl          (0),
		.gen3_coeff_10_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_10_nxtber_more_hwtcl          ("g3_coeff_10_nxtber_more"),
		.gen3_coeff_10_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_10_nxtber_less_hwtcl          ("g3_coeff_10_nxtber_less"),
		.gen3_coeff_10_reqber_hwtcl               (0),
		.gen3_coeff_10_ber_meas_hwtcl             (0),
		.gen3_coeff_11_hwtcl                      (0),
		.gen3_coeff_11_sel_hwtcl                  ("preset_11"),
		.gen3_coeff_11_preset_hint_hwtcl          (0),
		.gen3_coeff_11_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_11_nxtber_more_hwtcl          ("g3_coeff_11_nxtber_more"),
		.gen3_coeff_11_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_11_nxtber_less_hwtcl          ("g3_coeff_11_nxtber_less"),
		.gen3_coeff_11_reqber_hwtcl               (0),
		.gen3_coeff_11_ber_meas_hwtcl             (0),
		.gen3_coeff_12_hwtcl                      (0),
		.gen3_coeff_12_sel_hwtcl                  ("preset_12"),
		.gen3_coeff_12_preset_hint_hwtcl          (0),
		.gen3_coeff_12_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_12_nxtber_more_hwtcl          ("g3_coeff_12_nxtber_more"),
		.gen3_coeff_12_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_12_nxtber_less_hwtcl          ("g3_coeff_12_nxtber_less"),
		.gen3_coeff_12_reqber_hwtcl               (0),
		.gen3_coeff_12_ber_meas_hwtcl             (0),
		.gen3_coeff_13_hwtcl                      (0),
		.gen3_coeff_13_sel_hwtcl                  ("preset_13"),
		.gen3_coeff_13_preset_hint_hwtcl          (0),
		.gen3_coeff_13_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_13_nxtber_more_hwtcl          ("g3_coeff_13_nxtber_more"),
		.gen3_coeff_13_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_13_nxtber_less_hwtcl          ("g3_coeff_13_nxtber_less"),
		.gen3_coeff_13_reqber_hwtcl               (0),
		.gen3_coeff_13_ber_meas_hwtcl             (0),
		.gen3_coeff_14_hwtcl                      (0),
		.gen3_coeff_14_sel_hwtcl                  ("preset_14"),
		.gen3_coeff_14_preset_hint_hwtcl          (0),
		.gen3_coeff_14_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_14_nxtber_more_hwtcl          ("g3_coeff_14_nxtber_more"),
		.gen3_coeff_14_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_14_nxtber_less_hwtcl          ("g3_coeff_14_nxtber_less"),
		.gen3_coeff_14_reqber_hwtcl               (0),
		.gen3_coeff_14_ber_meas_hwtcl             (0),
		.gen3_coeff_15_hwtcl                      (0),
		.gen3_coeff_15_sel_hwtcl                  ("preset_15"),
		.gen3_coeff_15_preset_hint_hwtcl          (0),
		.gen3_coeff_15_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_15_nxtber_more_hwtcl          ("g3_coeff_15_nxtber_more"),
		.gen3_coeff_15_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_15_nxtber_less_hwtcl          ("g3_coeff_15_nxtber_less"),
		.gen3_coeff_15_reqber_hwtcl               (0),
		.gen3_coeff_15_ber_meas_hwtcl             (0),
		.gen3_coeff_16_hwtcl                      (0),
		.gen3_coeff_16_sel_hwtcl                  ("preset_16"),
		.gen3_coeff_16_preset_hint_hwtcl          (0),
		.gen3_coeff_16_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_16_nxtber_more_hwtcl          ("g3_coeff_16_nxtber_more"),
		.gen3_coeff_16_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_16_nxtber_less_hwtcl          ("g3_coeff_16_nxtber_less"),
		.gen3_coeff_16_reqber_hwtcl               (0),
		.gen3_coeff_16_ber_meas_hwtcl             (0),
		.gen3_coeff_17_hwtcl                      (0),
		.gen3_coeff_17_sel_hwtcl                  ("preset_17"),
		.gen3_coeff_17_preset_hint_hwtcl          (0),
		.gen3_coeff_17_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_17_nxtber_more_hwtcl          ("g3_coeff_17_nxtber_more"),
		.gen3_coeff_17_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_17_nxtber_less_hwtcl          ("g3_coeff_17_nxtber_less"),
		.gen3_coeff_17_reqber_hwtcl               (0),
		.gen3_coeff_17_ber_meas_hwtcl             (0),
		.gen3_coeff_18_hwtcl                      (0),
		.gen3_coeff_18_sel_hwtcl                  ("preset_18"),
		.gen3_coeff_18_preset_hint_hwtcl          (0),
		.gen3_coeff_18_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_18_nxtber_more_hwtcl          ("g3_coeff_18_nxtber_more"),
		.gen3_coeff_18_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_18_nxtber_less_hwtcl          ("g3_coeff_18_nxtber_less"),
		.gen3_coeff_18_reqber_hwtcl               (0),
		.gen3_coeff_18_ber_meas_hwtcl             (0),
		.gen3_coeff_19_hwtcl                      (0),
		.gen3_coeff_19_sel_hwtcl                  ("preset_19"),
		.gen3_coeff_19_preset_hint_hwtcl          (0),
		.gen3_coeff_19_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_19_nxtber_more_hwtcl          ("g3_coeff_19_nxtber_more"),
		.gen3_coeff_19_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_19_nxtber_less_hwtcl          ("g3_coeff_19_nxtber_less"),
		.gen3_coeff_19_reqber_hwtcl               (0),
		.gen3_coeff_19_ber_meas_hwtcl             (0),
		.gen3_coeff_20_hwtcl                      (0),
		.gen3_coeff_20_sel_hwtcl                  ("preset_20"),
		.gen3_coeff_20_preset_hint_hwtcl          (0),
		.gen3_coeff_20_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_20_nxtber_more_hwtcl          ("g3_coeff_20_nxtber_more"),
		.gen3_coeff_20_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_20_nxtber_less_hwtcl          ("g3_coeff_20_nxtber_less"),
		.gen3_coeff_20_reqber_hwtcl               (0),
		.gen3_coeff_20_ber_meas_hwtcl             (0),
		.gen3_coeff_21_hwtcl                      (0),
		.gen3_coeff_21_sel_hwtcl                  ("preset_21"),
		.gen3_coeff_21_preset_hint_hwtcl          (0),
		.gen3_coeff_21_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_21_nxtber_more_hwtcl          ("g3_coeff_21_nxtber_more"),
		.gen3_coeff_21_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_21_nxtber_less_hwtcl          ("g3_coeff_21_nxtber_less"),
		.gen3_coeff_21_reqber_hwtcl               (0),
		.gen3_coeff_21_ber_meas_hwtcl             (0),
		.gen3_coeff_22_hwtcl                      (0),
		.gen3_coeff_22_sel_hwtcl                  ("preset_22"),
		.gen3_coeff_22_preset_hint_hwtcl          (0),
		.gen3_coeff_22_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_22_nxtber_more_hwtcl          ("g3_coeff_22_nxtber_more"),
		.gen3_coeff_22_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_22_nxtber_less_hwtcl          ("g3_coeff_22_nxtber_less"),
		.gen3_coeff_22_reqber_hwtcl               (0),
		.gen3_coeff_22_ber_meas_hwtcl             (0),
		.gen3_coeff_23_hwtcl                      (0),
		.gen3_coeff_23_sel_hwtcl                  ("preset_23"),
		.gen3_coeff_23_preset_hint_hwtcl          (0),
		.gen3_coeff_23_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_23_nxtber_more_hwtcl          ("g3_coeff_23_nxtber_more"),
		.gen3_coeff_23_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_23_nxtber_less_hwtcl          ("g3_coeff_23_nxtber_less"),
		.gen3_coeff_23_reqber_hwtcl               (0),
		.gen3_coeff_23_ber_meas_hwtcl             (0),
		.gen3_coeff_24_hwtcl                      (0),
		.gen3_coeff_24_sel_hwtcl                  ("preset_24"),
		.gen3_coeff_24_preset_hint_hwtcl          (0),
		.gen3_coeff_24_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_24_nxtber_more_hwtcl          ("g3_coeff_24_nxtber_more"),
		.gen3_coeff_24_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_24_nxtber_less_hwtcl          ("g3_coeff_24_nxtber_less"),
		.gen3_coeff_24_reqber_hwtcl               (0),
		.gen3_coeff_24_ber_meas_hwtcl             (0),
		.hwtcl_override_g3txcoef                  (0),
		.gen3_preset_coeff_1_hwtcl                (0),
		.gen3_preset_coeff_2_hwtcl                (0),
		.gen3_preset_coeff_3_hwtcl                (0),
		.gen3_preset_coeff_4_hwtcl                (0),
		.gen3_preset_coeff_5_hwtcl                (0),
		.gen3_preset_coeff_6_hwtcl                (0),
		.gen3_preset_coeff_7_hwtcl                (0),
		.gen3_preset_coeff_8_hwtcl                (0),
		.gen3_preset_coeff_9_hwtcl                (0),
		.gen3_preset_coeff_10_hwtcl               (0),
		.gen3_preset_coeff_11_hwtcl               (0),
		.gen3_low_freq_hwtcl                      (0),
		.full_swing_hwtcl                         (35),
		.gen3_full_swing_hwtcl                    (35),
		.use_atx_pll_hwtcl                        (0),
		.low_latency_mode_hwtcl                   (0)
	) dut (
		.npor                   (pcie_rstn_npor),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //               npor.npor
		.pin_perst              (pcie_rstn_pin_perst),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .pin_perst
		.lmi_addr               (apps_lmi_lmi_addr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                lmi.lmi_addr
		.lmi_din                (apps_lmi_lmi_din),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .lmi_din
		.lmi_rden               (apps_lmi_lmi_rden),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .lmi_rden
		.lmi_wren               (apps_lmi_lmi_wren),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .lmi_wren
		.lmi_ack                (dut_lmi_lmi_ack),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .lmi_ack
		.lmi_dout               (dut_lmi_lmi_dout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .lmi_dout
		.hpg_ctrler             (apps_config_tl_hpg_ctrler),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //          config_tl.hpg_ctrler
		.tl_cfg_add             (dut_config_tl_tl_cfg_add),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .tl_cfg_add
		.tl_cfg_ctl             (dut_config_tl_tl_cfg_ctl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .tl_cfg_ctl
		.tl_cfg_sts             (dut_config_tl_tl_cfg_sts),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .tl_cfg_sts
		.cpl_err                (apps_config_tl_cpl_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .cpl_err
		.cpl_pending            (apps_config_tl_cpl_pending),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .cpl_pending
		.pm_auxpwr              (apps_power_mngt_pm_auxpwr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //         power_mngt.pm_auxpwr
		.pm_data                (apps_power_mngt_pm_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .pm_data
		.pme_to_cr              (apps_power_mngt_pme_to_cr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .pme_to_cr
		.pm_event               (apps_power_mngt_pm_event),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .pm_event
		.pme_to_sr              (dut_power_mngt_pme_to_sr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .pme_to_sr
		.rx_st_sop              (dut_rx_st_startofpacket),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //              rx_st.startofpacket
		.rx_st_eop              (dut_rx_st_endofpacket),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                   .endofpacket
		.rx_st_err              (dut_rx_st_error),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .error
		.rx_st_valid            (dut_rx_st_valid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .valid
		.rx_st_empty            (dut_rx_st_empty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .empty
		.rx_st_ready            (dut_rx_st_ready),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .ready
		.rx_st_data             (dut_rx_st_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .data
		.rx_st_bar              (dut_rx_bar_be_rx_st_bar),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //          rx_bar_be.rx_st_bar
		.rx_st_be               (dut_rx_bar_be_rx_st_be),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .rx_st_be
		.rx_st_mask             (apps_rx_bar_be_rx_st_mask),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rx_st_mask
		.tx_st_sop              (apps_tx_st_startofpacket),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //              tx_st.startofpacket
		.tx_st_eop              (apps_tx_st_endofpacket),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .endofpacket
		.tx_st_err              (apps_tx_st_error),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .error
		.tx_st_valid            (apps_tx_st_valid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .valid
		.tx_st_empty            (apps_tx_st_empty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .empty
		.tx_st_ready            (apps_tx_st_ready),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .ready
		.tx_st_data             (apps_tx_st_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .data
		.tx_cred_datafccp       (dut_tx_cred_tx_cred_datafccp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //            tx_cred.tx_cred_datafccp
		.tx_cred_datafcnp       (dut_tx_cred_tx_cred_datafcnp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //                   .tx_cred_datafcnp
		.tx_cred_datafcp        (dut_tx_cred_tx_cred_datafcp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .tx_cred_datafcp
		.tx_cred_fchipcons      (dut_tx_cred_tx_cred_fchipcons),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .tx_cred_fchipcons
		.tx_cred_fcinfinite     (dut_tx_cred_tx_cred_fcinfinite),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .tx_cred_fcinfinite
		.tx_cred_hdrfccp        (dut_tx_cred_tx_cred_hdrfccp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .tx_cred_hdrfccp
		.tx_cred_hdrfcnp        (dut_tx_cred_tx_cred_hdrfcnp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .tx_cred_hdrfcnp
		.tx_cred_hdrfcp         (dut_tx_cred_tx_cred_hdrfcp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .tx_cred_hdrfcp
		.pld_clk                (apps_pld_clk_hip_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //            pld_clk.clk
		.coreclkout_hip         (dut_coreclkout_hip_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //     coreclkout_hip.clk
		.refclk                 (refclk_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //             refclk.clk
		.reset_status           (dut_hip_rst_reset_status),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //            hip_rst.reset_status
		.serdes_pll_locked      (dut_hip_rst_serdes_pll_locked),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .serdes_pll_locked
		.pld_clk_inuse          (dut_hip_rst_pld_clk_inuse),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .pld_clk_inuse
		.pld_core_ready         (apps_hip_rst_pld_core_ready),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .pld_core_ready
		.testin_zero            (dut_hip_rst_testin_zero),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .testin_zero
		.reconfig_to_xcvr       (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr     (dut_reconfig_from_xcvr_reconfig_from_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       // reconfig_from_xcvr.reconfig_from_xcvr
		.rx_in0                 (hip_serial_rx_in0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //         hip_serial.rx_in0
		.rx_in1                 (hip_serial_rx_in1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rx_in1
		.rx_in2                 (hip_serial_rx_in2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rx_in2
		.rx_in3                 (hip_serial_rx_in3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rx_in3
		.rx_in4                 (hip_serial_rx_in4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rx_in4
		.rx_in5                 (hip_serial_rx_in5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rx_in5
		.rx_in6                 (hip_serial_rx_in6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rx_in6
		.rx_in7                 (hip_serial_rx_in7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rx_in7
		.tx_out0                (hip_serial_tx_out0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_out0
		.tx_out1                (hip_serial_tx_out1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_out1
		.tx_out2                (hip_serial_tx_out2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_out2
		.tx_out3                (hip_serial_tx_out3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_out3
		.tx_out4                (hip_serial_tx_out4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_out4
		.tx_out5                (hip_serial_tx_out5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_out5
		.tx_out6                (hip_serial_tx_out6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_out6
		.tx_out7                (hip_serial_tx_out7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_out7
		.sim_pipe_pclk_in       (hip_pipe_sim_pipe_pclk_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //           hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate          (hip_pipe_sim_pipe_rate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .sim_pipe_rate
		.sim_ltssmstate         (hip_pipe_sim_ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .sim_ltssmstate
		.eidleinfersel0         (hip_pipe_eidleinfersel0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel0
		.eidleinfersel1         (hip_pipe_eidleinfersel1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel1
		.eidleinfersel2         (hip_pipe_eidleinfersel2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel2
		.eidleinfersel3         (hip_pipe_eidleinfersel3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel3
		.eidleinfersel4         (hip_pipe_eidleinfersel4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel4
		.eidleinfersel5         (hip_pipe_eidleinfersel5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel5
		.eidleinfersel6         (hip_pipe_eidleinfersel6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel6
		.eidleinfersel7         (hip_pipe_eidleinfersel7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .eidleinfersel7
		.powerdown0             (hip_pipe_powerdown0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown0
		.powerdown1             (hip_pipe_powerdown1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown1
		.powerdown2             (hip_pipe_powerdown2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown2
		.powerdown3             (hip_pipe_powerdown3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown3
		.powerdown4             (hip_pipe_powerdown4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown4
		.powerdown5             (hip_pipe_powerdown5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown5
		.powerdown6             (hip_pipe_powerdown6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown6
		.powerdown7             (hip_pipe_powerdown7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .powerdown7
		.rxpolarity0            (hip_pipe_rxpolarity0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity0
		.rxpolarity1            (hip_pipe_rxpolarity1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity1
		.rxpolarity2            (hip_pipe_rxpolarity2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity2
		.rxpolarity3            (hip_pipe_rxpolarity3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity3
		.rxpolarity4            (hip_pipe_rxpolarity4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity4
		.rxpolarity5            (hip_pipe_rxpolarity5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity5
		.rxpolarity6            (hip_pipe_rxpolarity6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity6
		.rxpolarity7            (hip_pipe_rxpolarity7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxpolarity7
		.txcompl0               (hip_pipe_txcompl0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl0
		.txcompl1               (hip_pipe_txcompl1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl1
		.txcompl2               (hip_pipe_txcompl2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl2
		.txcompl3               (hip_pipe_txcompl3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl3
		.txcompl4               (hip_pipe_txcompl4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl4
		.txcompl5               (hip_pipe_txcompl5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl5
		.txcompl6               (hip_pipe_txcompl6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl6
		.txcompl7               (hip_pipe_txcompl7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txcompl7
		.txdata0                (hip_pipe_txdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata0
		.txdata1                (hip_pipe_txdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata1
		.txdata2                (hip_pipe_txdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata2
		.txdata3                (hip_pipe_txdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata3
		.txdata4                (hip_pipe_txdata4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata4
		.txdata5                (hip_pipe_txdata5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata5
		.txdata6                (hip_pipe_txdata6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata6
		.txdata7                (hip_pipe_txdata7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .txdata7
		.txdatak0               (hip_pipe_txdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak0
		.txdatak1               (hip_pipe_txdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak1
		.txdatak2               (hip_pipe_txdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak2
		.txdatak3               (hip_pipe_txdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak3
		.txdatak4               (hip_pipe_txdatak4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak4
		.txdatak5               (hip_pipe_txdatak5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak5
		.txdatak6               (hip_pipe_txdatak6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak6
		.txdatak7               (hip_pipe_txdatak7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txdatak7
		.txdetectrx0            (hip_pipe_txdetectrx0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx0
		.txdetectrx1            (hip_pipe_txdetectrx1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx1
		.txdetectrx2            (hip_pipe_txdetectrx2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx2
		.txdetectrx3            (hip_pipe_txdetectrx3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx3
		.txdetectrx4            (hip_pipe_txdetectrx4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx4
		.txdetectrx5            (hip_pipe_txdetectrx5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx5
		.txdetectrx6            (hip_pipe_txdetectrx6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx6
		.txdetectrx7            (hip_pipe_txdetectrx7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txdetectrx7
		.txelecidle0            (hip_pipe_txelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle0
		.txelecidle1            (hip_pipe_txelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle1
		.txelecidle2            (hip_pipe_txelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle2
		.txelecidle3            (hip_pipe_txelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle3
		.txelecidle4            (hip_pipe_txelecidle4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle4
		.txelecidle5            (hip_pipe_txelecidle5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle5
		.txelecidle6            (hip_pipe_txelecidle6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle6
		.txelecidle7            (hip_pipe_txelecidle7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .txelecidle7
		.txdeemph0              (hip_pipe_txdeemph0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph0
		.txdeemph1              (hip_pipe_txdeemph1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph1
		.txdeemph2              (hip_pipe_txdeemph2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph2
		.txdeemph3              (hip_pipe_txdeemph3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph3
		.txdeemph4              (hip_pipe_txdeemph4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph4
		.txdeemph5              (hip_pipe_txdeemph5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph5
		.txdeemph6              (hip_pipe_txdeemph6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph6
		.txdeemph7              (hip_pipe_txdeemph7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txdeemph7
		.txmargin0              (hip_pipe_txmargin0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin0
		.txmargin1              (hip_pipe_txmargin1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin1
		.txmargin2              (hip_pipe_txmargin2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin2
		.txmargin3              (hip_pipe_txmargin3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin3
		.txmargin4              (hip_pipe_txmargin4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin4
		.txmargin5              (hip_pipe_txmargin5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin5
		.txmargin6              (hip_pipe_txmargin6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin6
		.txmargin7              (hip_pipe_txmargin7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .txmargin7
		.txswing0               (hip_pipe_txswing0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing0
		.txswing1               (hip_pipe_txswing1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing1
		.txswing2               (hip_pipe_txswing2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing2
		.txswing3               (hip_pipe_txswing3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing3
		.txswing4               (hip_pipe_txswing4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing4
		.txswing5               (hip_pipe_txswing5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing5
		.txswing6               (hip_pipe_txswing6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing6
		.txswing7               (hip_pipe_txswing7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .txswing7
		.phystatus0             (hip_pipe_phystatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus0
		.phystatus1             (hip_pipe_phystatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus1
		.phystatus2             (hip_pipe_phystatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus2
		.phystatus3             (hip_pipe_phystatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus3
		.phystatus4             (hip_pipe_phystatus4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus4
		.phystatus5             (hip_pipe_phystatus5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus5
		.phystatus6             (hip_pipe_phystatus6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus6
		.phystatus7             (hip_pipe_phystatus7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .phystatus7
		.rxdata0                (hip_pipe_rxdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata0
		.rxdata1                (hip_pipe_rxdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata1
		.rxdata2                (hip_pipe_rxdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata2
		.rxdata3                (hip_pipe_rxdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata3
		.rxdata4                (hip_pipe_rxdata4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata4
		.rxdata5                (hip_pipe_rxdata5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata5
		.rxdata6                (hip_pipe_rxdata6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata6
		.rxdata7                (hip_pipe_rxdata7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .rxdata7
		.rxdatak0               (hip_pipe_rxdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak0
		.rxdatak1               (hip_pipe_rxdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak1
		.rxdatak2               (hip_pipe_rxdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak2
		.rxdatak3               (hip_pipe_rxdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak3
		.rxdatak4               (hip_pipe_rxdatak4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak4
		.rxdatak5               (hip_pipe_rxdatak5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak5
		.rxdatak6               (hip_pipe_rxdatak6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak6
		.rxdatak7               (hip_pipe_rxdatak7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxdatak7
		.rxelecidle0            (hip_pipe_rxelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle0
		.rxelecidle1            (hip_pipe_rxelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle1
		.rxelecidle2            (hip_pipe_rxelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle2
		.rxelecidle3            (hip_pipe_rxelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle3
		.rxelecidle4            (hip_pipe_rxelecidle4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle4
		.rxelecidle5            (hip_pipe_rxelecidle5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle5
		.rxelecidle6            (hip_pipe_rxelecidle6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle6
		.rxelecidle7            (hip_pipe_rxelecidle7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .rxelecidle7
		.rxstatus0              (hip_pipe_rxstatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus0
		.rxstatus1              (hip_pipe_rxstatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus1
		.rxstatus2              (hip_pipe_rxstatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus2
		.rxstatus3              (hip_pipe_rxstatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus3
		.rxstatus4              (hip_pipe_rxstatus4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus4
		.rxstatus5              (hip_pipe_rxstatus5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus5
		.rxstatus6              (hip_pipe_rxstatus6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus6
		.rxstatus7              (hip_pipe_rxstatus7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .rxstatus7
		.rxvalid0               (hip_pipe_rxvalid0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid0
		.rxvalid1               (hip_pipe_rxvalid1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid1
		.rxvalid2               (hip_pipe_rxvalid2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid2
		.rxvalid3               (hip_pipe_rxvalid3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid3
		.rxvalid4               (hip_pipe_rxvalid4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid4
		.rxvalid5               (hip_pipe_rxvalid5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid5
		.rxvalid6               (hip_pipe_rxvalid6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid6
		.rxvalid7               (hip_pipe_rxvalid7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .rxvalid7
		.app_int_sts            (apps_int_msi_app_int_sts),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //            int_msi.app_int_sts
		.app_msi_num            (apps_int_msi_app_msi_num),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .app_msi_num
		.app_msi_req            (apps_int_msi_app_msi_req),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .app_msi_req
		.app_msi_tc             (apps_int_msi_app_msi_tc),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .app_msi_tc
		.app_int_ack            (dut_int_msi_app_int_ack),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .app_int_ack
		.app_msi_ack            (dut_int_msi_app_msi_ack),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .app_msi_ack
		.test_in                (hip_ctrl_test_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           hip_ctrl.test_in
		.simu_mode_pipe         (hip_ctrl_simu_mode_pipe),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .simu_mode_pipe
		.derr_cor_ext_rcv       (dut_hip_status_derr_cor_ext_rcv),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //         hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl       (dut_hip_status_derr_cor_ext_rpl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .derr_cor_ext_rpl
		.derr_rpl               (dut_hip_status_derr_rpl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .derr_rpl
		.dlup                   (dut_hip_status_dlup),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             //                   .dlup
		.dlup_exit              (dut_hip_status_dlup_exit),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .dlup_exit
		.ev128ns                (dut_hip_status_ev128ns),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .ev128ns
		.ev1us                  (dut_hip_status_ev1us),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .ev1us
		.hotrst_exit            (dut_hip_status_hotrst_exit),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .hotrst_exit
		.int_status             (dut_hip_status_int_status),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .int_status
		.l2_exit                (dut_hip_status_l2_exit),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .l2_exit
		.lane_act               (dut_hip_status_lane_act),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .lane_act
		.ltssmstate             (dut_hip_status_ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .ltssmstate
		.rx_par_err             (dut_hip_status_rx_par_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rx_par_err
		.tx_par_err             (dut_hip_status_tx_par_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .tx_par_err
		.cfg_par_err            (dut_hip_status_cfg_par_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .cfg_par_err
		.ko_cpl_spc_header      (dut_hip_status_ko_cpl_spc_header),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .ko_cpl_spc_header
		.ko_cpl_spc_data        (dut_hip_status_ko_cpl_spc_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .ko_cpl_spc_data
		.currentspeed           (dut_hip_currentspeed_currentspeed),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //   hip_currentspeed.currentspeed
		.rx_st_parity           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.tx_st_parity           (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.sim_pipe_pclk_out      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.rxdataskip0            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip1            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip2            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip3            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip4            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip5            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip6            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip7            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst0               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst1               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst2               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst3               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst4               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst5               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst6               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst7               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxsynchd0              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd1              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd2              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd3              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd4              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd5              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd6              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd7              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxfreqlocked0          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked1          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked2          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked3          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked4          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked5          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked6          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked7          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.currentcoeff0          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff1          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff2          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff3          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff4          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff5          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff6          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff7          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset0       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset1       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset2       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset3       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset4       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset5       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset6       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset7       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd0              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd1              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd2              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd3              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst0               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst1               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst2               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst3               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst4               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst5               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst6               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst7               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.aer_msi_num            (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.pex_msi_num            (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.serr_out               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.hip_reconfig_clk       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_rst_n     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_address   (10'b0000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //        (terminated)
		.hip_reconfig_read      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_write     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_writedata (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_byte_en   (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.ser_shift_load         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.interface_sel          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_link2csr         (13'b0000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //        (terminated)
		.cfgbp_comclk_reg       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_extsy_reg        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_max_pload        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
		.cfgbp_tx_ecrcgen       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_rx_ecrchk        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_secbus           (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //        (terminated)
		.cfgbp_linkcsr_bit0     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_tx_req_pm        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_tx_typ_pm        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
		.cfgbp_req_phypm        (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
		.cfgbp_req_phycfg       (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
		.cfgbp_vc0_tcmap_pld    (7'b0000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //        (terminated)
		.cfgbp_inh_dllp         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_inh_tx_tlp       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_req_wake         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_link3_ctl        (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.cseb_rddata            (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cseb_rdresponse        (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.cseb_waitrequest       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cseb_wrresponse        (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.cseb_wrresp_valid      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cseb_rddata_parity     (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
		.reservedin             (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.tlbfm_in               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.tlbfm_out              (1001'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.rxfc_cplbuf_ovf        ()                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //        (terminated)
	);

	altpcied_sv_hwtcl #(
		.device_family_hwtcl              ("Stratix V"),
		.lane_mask_hwtcl                  ("x8"),
		.gen123_lane_rate_mode_hwtcl      ("Gen1 (2.5 Gbps)"),
		.pld_clockrate_hwtcl              (125000000),
		.port_type_hwtcl                  ("Native endpoint"),
		.ast_width_hwtcl                  ("Avalon-ST 128-bit"),
		.extend_tag_field_hwtcl           (32),
		.max_payload_size_hwtcl           (256),
		.num_of_func_hwtcl                (1),
		.multiple_packets_per_cycle_hwtcl (0),
		.port_width_be_hwtcl              (16),
		.port_width_data_hwtcl            (128),
		.avalon_waddr_hwltcl              (12),
		.check_bus_master_ena_hwtcl       (1),
		.check_rx_buffer_cpl_hwtcl        (1),
		.use_crc_forwarding_hwtcl         (0)
	) apps (
		.coreclkout_hip       (dut_coreclkout_hip_clk),                   // coreclkout_hip.clk
		.pld_clk_hip          (apps_pld_clk_hip_clk),                     //    pld_clk_hip.clk
		.rx_st_sop            (dut_rx_st_startofpacket),                  //          rx_st.startofpacket
		.rx_st_eop            (dut_rx_st_endofpacket),                    //               .endofpacket
		.rx_st_err            (dut_rx_st_error),                          //               .error
		.rx_st_valid          (dut_rx_st_valid),                          //               .valid
		.rx_st_empty          (dut_rx_st_empty),                          //               .empty
		.rx_st_ready          (dut_rx_st_ready),                          //               .ready
		.rx_st_data           (dut_rx_st_data),                           //               .data
		.rx_st_bar            (dut_rx_bar_be_rx_st_bar),                  //      rx_bar_be.rx_st_bar
		.rx_st_be             (dut_rx_bar_be_rx_st_be),                   //               .rx_st_be
		.rx_st_mask           (apps_rx_bar_be_rx_st_mask),                //               .rx_st_mask
		.tx_st_sop            (apps_tx_st_startofpacket),                 //          tx_st.startofpacket
		.tx_st_eop            (apps_tx_st_endofpacket),                   //               .endofpacket
		.tx_st_err            (apps_tx_st_error),                         //               .error
		.tx_st_valid          (apps_tx_st_valid),                         //               .valid
		.tx_st_empty          (apps_tx_st_empty),                         //               .empty
		.tx_st_ready          (apps_tx_st_ready),                         //               .ready
		.tx_st_data           (apps_tx_st_data),                          //               .data
		.tx_cred_datafccp     (dut_tx_cred_tx_cred_datafccp),             //        tx_cred.tx_cred_datafccp
		.tx_cred_datafcnp     (dut_tx_cred_tx_cred_datafcnp),             //               .tx_cred_datafcnp
		.tx_cred_datafcp      (dut_tx_cred_tx_cred_datafcp),              //               .tx_cred_datafcp
		.tx_cred_fchipcons    (dut_tx_cred_tx_cred_fchipcons),            //               .tx_cred_fchipcons
		.tx_cred_fcinfinite   (dut_tx_cred_tx_cred_fcinfinite),           //               .tx_cred_fcinfinite
		.tx_cred_hdrfccp      (dut_tx_cred_tx_cred_hdrfccp),              //               .tx_cred_hdrfccp
		.tx_cred_hdrfcnp      (dut_tx_cred_tx_cred_hdrfcnp),              //               .tx_cred_hdrfcnp
		.tx_cred_hdrfcp       (dut_tx_cred_tx_cred_hdrfcp),               //               .tx_cred_hdrfcp
		.reset_status         (dut_hip_rst_reset_status),                 //        hip_rst.reset_status
		.serdes_pll_locked    (dut_hip_rst_serdes_pll_locked),            //               .serdes_pll_locked
		.pld_clk_inuse        (dut_hip_rst_pld_clk_inuse),                //               .pld_clk_inuse
		.pld_core_ready       (apps_hip_rst_pld_core_ready),              //               .pld_core_ready
		.testin_zero          (dut_hip_rst_testin_zero),                  //               .testin_zero
		.app_int_sts          (apps_int_msi_app_int_sts),                 //        int_msi.app_int_sts
		.app_int_ack          (dut_int_msi_app_int_ack),                  //               .app_int_ack
		.app_msi_req          (apps_int_msi_app_msi_req),                 //               .app_msi_req
		.app_msi_tc           (apps_int_msi_app_msi_tc),                  //               .app_msi_tc
		.app_msi_ack          (dut_int_msi_app_msi_ack),                  //               .app_msi_ack
		.app_msi_num          (apps_int_msi_app_msi_num),                 //               .app_msi_num
		.derr_cor_ext_rcv     (dut_hip_status_derr_cor_ext_rcv),          //     hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl     (dut_hip_status_derr_cor_ext_rpl),          //               .derr_cor_ext_rpl
		.derr_rpl             (dut_hip_status_derr_rpl),                  //               .derr_rpl
		.dlup_exit            (dut_hip_status_dlup_exit),                 //               .dlup_exit
		.ev128ns              (dut_hip_status_ev128ns),                   //               .ev128ns
		.ev1us                (dut_hip_status_ev1us),                     //               .ev1us
		.hotrst_exit          (dut_hip_status_hotrst_exit),               //               .hotrst_exit
		.int_status           (dut_hip_status_int_status),                //               .int_status
		.l2_exit              (dut_hip_status_l2_exit),                   //               .l2_exit
		.lane_act             (dut_hip_status_lane_act),                  //               .lane_act
		.ltssmstate           (dut_hip_status_ltssmstate),                //               .ltssmstate
		.dlup                 (dut_hip_status_dlup),                      //               .dlup
		.rx_par_err           (dut_hip_status_rx_par_err),                //               .rx_par_err
		.tx_par_err           (dut_hip_status_tx_par_err),                //               .tx_par_err
		.cfg_par_err          (dut_hip_status_cfg_par_err),               //               .cfg_par_err
		.ko_cpl_spc_header    (dut_hip_status_ko_cpl_spc_header),         //               .ko_cpl_spc_header
		.ko_cpl_spc_data      (dut_hip_status_ko_cpl_spc_data),           //               .ko_cpl_spc_data
		.derr_cor_ext_rcv_drv (apps_hip_status_drv_derr_cor_ext_rcv_drv), // hip_status_drv.derr_cor_ext_rcv_drv
		.derr_cor_ext_rpl_drv (apps_hip_status_drv_derr_cor_ext_rpl_drv), //               .derr_cor_ext_rpl_drv
		.derr_rpl_drv         (apps_hip_status_drv_derr_rpl_drv),         //               .derr_rpl_drv
		.dlup_exit_drv        (apps_hip_status_drv_dlup_exit_drv),        //               .dlup_exit_drv
		.ev128ns_drv          (apps_hip_status_drv_ev128ns_drv),          //               .ev128ns_drv
		.ev1us_drv            (apps_hip_status_drv_ev1us_drv),            //               .ev1us_drv
		.hotrst_exit_drv      (apps_hip_status_drv_hotrst_exit_drv),      //               .hotrst_exit_drv
		.int_status_drv       (apps_hip_status_drv_int_status_drv),       //               .int_status_drv
		.l2_exit_drv          (apps_hip_status_drv_l2_exit_drv),          //               .l2_exit_drv
		.lane_act_drv         (apps_hip_status_drv_lane_act_drv),         //               .lane_act_drv
		.ltssmstate_drv       (apps_hip_status_drv_ltssmstate_drv),       //               .ltssmstate_drv
		.hpg_ctrler           (apps_config_tl_hpg_ctrler),                //      config_tl.hpg_ctrler
		.tl_cfg_ctl           (dut_config_tl_tl_cfg_ctl),                 //               .tl_cfg_ctl
		.cpl_err              (apps_config_tl_cpl_err),                   //               .cpl_err
		.tl_cfg_add           (dut_config_tl_tl_cfg_add),                 //               .tl_cfg_add
		.tl_cfg_sts           (dut_config_tl_tl_cfg_sts),                 //               .tl_cfg_sts
		.cpl_pending          (apps_config_tl_cpl_pending),               //               .cpl_pending
		.lmi_addr             (apps_lmi_lmi_addr),                        //            lmi.lmi_addr
		.lmi_din              (apps_lmi_lmi_din),                         //               .lmi_din
		.lmi_rden             (apps_lmi_lmi_rden),                        //               .lmi_rden
		.lmi_wren             (apps_lmi_lmi_wren),                        //               .lmi_wren
		.lmi_ack              (dut_lmi_lmi_ack),                          //               .lmi_ack
		.lmi_dout             (dut_lmi_lmi_dout),                         //               .lmi_dout
		.pm_auxpwr            (apps_power_mngt_pm_auxpwr),                //     power_mngt.pm_auxpwr
		.pm_data              (apps_power_mngt_pm_data),                  //               .pm_data
		.pme_to_cr            (apps_power_mngt_pme_to_cr),                //               .pme_to_cr
		.pm_event             (apps_power_mngt_pm_event),                 //               .pm_event
		.pme_to_sr            (dut_power_mngt_pme_to_sr),                 //               .pme_to_sr
		.rx_st_parity         (16'b0000000000000000),                     //    (terminated)
		.rx_bar_dec_func_num  (3'b000),                                   //    (terminated)
		.tx_st_parity         (),                                         //    (terminated)
		.tx_fifo_empty        (1'b1),                                     //    (terminated)
		.sim_pipe_pclk_out    (1'b0),                                     //    (terminated)
		.app_msi_func         (),                                         //    (terminated)
		.serr_out             (1'b0),                                     //    (terminated)
		.rxfc_cplbuf_ovf      (1'b0),                                     //    (terminated)
		.tl_cfg_ctl_wr        (1'b0),                                     //    (terminated)
		.tl_cfg_sts_wr        (1'b0),                                     //    (terminated)
		.cpl_err_func         (),                                         //    (terminated)
		.pm_event_func        ()                                          //    (terminated)
	);

	altpcie_reconfig_driver #(
		.gen123_lane_rate_mode_hwtcl   ("Gen1 (2.5 Gbps)"),
		.number_of_reconfig_interfaces (10)
	) pcie_reconfig_driver_0 (
		.reconfig_xcvr_clk         (clk_clk),                                          // reconfig_xcvr_clk.clk
		.reconfig_xcvr_rst         (rst_controller_reset_out_reset),                   // reconfig_xcvr_rst.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),     //     reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),        //                  .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),    //                  .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest), //                  .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),       //                  .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),   //                  .writedata
		.currentspeed              (dut_hip_currentspeed_currentspeed),                //  hip_currentspeed.currentspeed
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),  //     reconfig_busy.reconfig_busy
		.pld_clk                   (apps_pld_clk_hip_clk),                             //           pld_clk.clk
		.derr_cor_ext_rcv_drv      (apps_hip_status_drv_derr_cor_ext_rcv_drv),         //    hip_status_drv.derr_cor_ext_rcv_drv
		.derr_cor_ext_rpl_drv      (apps_hip_status_drv_derr_cor_ext_rpl_drv),         //                  .derr_cor_ext_rpl_drv
		.derr_rpl_drv              (apps_hip_status_drv_derr_rpl_drv),                 //                  .derr_rpl_drv
		.dlup_exit_drv             (apps_hip_status_drv_dlup_exit_drv),                //                  .dlup_exit_drv
		.ev128ns_drv               (apps_hip_status_drv_ev128ns_drv),                  //                  .ev128ns_drv
		.ev1us_drv                 (apps_hip_status_drv_ev1us_drv),                    //                  .ev1us_drv
		.hotrst_exit_drv           (apps_hip_status_drv_hotrst_exit_drv),              //                  .hotrst_exit_drv
		.int_status_drv            (apps_hip_status_drv_int_status_drv),               //                  .int_status_drv
		.l2_exit_drv               (apps_hip_status_drv_l2_exit_drv),                  //                  .l2_exit_drv
		.lane_act_drv              (apps_hip_status_drv_lane_act_drv),                 //                  .lane_act_drv
		.ltssmstate_drv            (apps_hip_status_drv_ltssmstate_drv)                //                  .ltssmstate_drv
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (10),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_analog                 (0),
		.enable_eyemon                 (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) alt_xcvr_reconfig_0 (
		.reconfig_busy             (alt_xcvr_reconfig_0_reconfig_busy_reconfig_busy),       //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_clk),                                               //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                        //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (pcie_reconfig_driver_0_reconfig_mgmt_address),          //      reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_reconfig_driver_0_reconfig_mgmt_read),             //                   .read
		.reconfig_mgmt_readdata    (pcie_reconfig_driver_0_reconfig_mgmt_readdata),         //                   .readdata
		.reconfig_mgmt_waitrequest (pcie_reconfig_driver_0_reconfig_mgmt_waitrequest),      //                   .waitrequest
		.reconfig_mgmt_write       (pcie_reconfig_driver_0_reconfig_mgmt_write),            //                   .write
		.reconfig_mgmt_writedata   (pcie_reconfig_driver_0_reconfig_mgmt_writedata),        //                   .writedata
		.reconfig_to_xcvr          (alt_xcvr_reconfig_0_reconfig_to_xcvr_reconfig_to_xcvr), //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (dut_reconfig_from_xcvr_reconfig_from_xcvr),             // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                      //        (terminated)
		.rx_cal_busy               (),                                                      //        (terminated)
		.cal_busy_in               (1'b0),                                                  //        (terminated)
		.reconfig_mif_address      (),                                                      //        (terminated)
		.reconfig_mif_read         (),                                                      //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                  //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                   //        (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
